library ieee;
use ieee.std_logic_1164.all;

entity LED_Blink is
end LED_Blink;

architecture RTL of LED_Blink is
begin
end architecture RTL;